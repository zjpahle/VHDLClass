library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity counter5bit_test is
end counter5bit_test;

architecture test of counter5bit_test is
--Signals Declarations--
	signal in1, rst	: std_logic;
	signal clk	: std_logic := '0';
	signal countOut	: std_logic_vector (4 downto 0);

--Component Instantiation--
	component counter5bit is
	port	(
		in1    		: in std_logic;
		rst    		: in std_logic;
		clk    		: in std_logic;
		countOut	: out std_logic_vector (4 downto 0)
		);

	end component counter5bit;

	begin counter5bit1 : counter5bit
	port map(
		in1		=> in1,
		rst		=> rst,
		clk		=> clk,
		countOut	=> countOut
		);

--Begin Testing--
	clk <= NOT clk after 1 ns;
	process begin
		in1 <= '0';
		rst <= '1';
		wait for 1 ns;
		rst <= '0';
		in1 <= '1';
		wait for 10 ns;
		in1 <= '0';
		wait for 2 ns;
		rst <= '1';
		wait for 1 ns;
	end process;

end architecture test;
