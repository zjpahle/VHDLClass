library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity memory8bit is
port	(
	rwsel, clk 	: in    std_logic;
	addr 		: in    std_logic_vector (7 downto 0);
	data    	: inout std_logic_vector (7 downto 0)
	);
end memory8bit;

architecture behavioral of memory8bit is
	type mem is array (natural range <>, natural range <>) of std_logic;
	constant memsize : integer := 2**addr'length;
	signal memory : mem (0 TO memsize-1, data'RANGE) :=  (others =>"00000000");
begin
	process (clk) begin
	if rising_edge(clk) then
		if (rwsel = '1') then
			for i in data'range loop
				data(i) <= memory(conv_integer(addr),i);
			end loop;
		else
			for i in data'range loop
				memory(conv_integer(addr),i) <= data(i);
			end loop;
		end if;
	end if;
	end process;
end behavioral;